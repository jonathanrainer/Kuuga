module load_store_unit(

    );
endmodule